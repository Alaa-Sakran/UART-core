`ifndef UART_HEADER_VH
`define UART_HEADER_VH
`include "AXI_UART_TX.v"
`include "clock_divider.v"
`include "fifo.v" 
`include "AXI_UART_RX.v"
`endif     
